module userInput();

// will be a counter from 0 - 12
/*
	0: null
	1:0
	2:1
	3:2
	...
	9:8
	10:9
	11:+
	12:-
	13:=
*/


endmodule
