module Lab6();

endmodule
