module pixelOutput();


/*
		// starting the vga output
		if (start == 1)
			startCount = startCount + 1;
		
		if (startCount == 10)
			begin	
				startCount = 0;
				vgaCount
*/

endmodule
