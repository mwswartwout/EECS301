module Lab4();

endmodule